module fivetothree_two_decoder_isd(d,a,enbl);
input [4:0]a;
input enbl;
output reg [31:0]d;
always @(a) 
  begin
    if(enbl==1)
      begin
        d[0] = !a[0] & !a[1] & !a[2] & !a[3] & !a[4];
        d[1] = a[0] & !a[1] & !a[2] & !a[3] & !a[4]; 
        d[2] = !a[0] & a[1] & !a[2] & !a[3] & !a[4];
        d[3] = a[0] & a[1] & !a[2] & !a[3] & !a[4];
        d[4] = !a[0] & !a[1] & a[2] & !a[3] & !a[4];
        d[5] = a[0] & !a[1] & a[2] & !a[3] & !a[4];
        d[6] = !a[0] & a[1] & a[2] & !a[3] & !a[4];
        d[7] = a[0] & a[1] & a[2] & !a[3] & !a[4];
        d[8] = !a[0] & !a[1] & !a[2] & a[3] & !a[4];
        d[9] = a[0] & !a[1] & !a[2] & a[3] & !a[4];
        d[10] = !a[0] & a[1] & !a[2] & a[3] & !a[4];
        d[11] = a[0] & a[1] & !a[2] & a[3] & !a[4]; 
        d[12] = !a[0] & !a[1] & a[2] & a[3] & !a[4];
        d[13] = a[0] & !a[1] & a[2] & a[3] & !a[4];
        d[14] = !a[0] & a[1] & a[2] & a[3] & !a[4];
        d[15] = a[0] & a[1] & a[2] & a[3] & !a[4];
        d[16] = !a[0] & !a[1] & !a[2] & !a[3] & a[4];
        d[17] = a[0] & !a[1] & !a[2] & !a[3] & a[4]; 
        d[18] = !a[0] & a[1] & !a[2] & !a[3] & a[4];
        d[19] = a[0] & a[1] & !a[2] & !a[3] & a[4];
        d[20] = !a[0] & !a[1] & a[2] & !a[3] & a[4];
        d[21] = a[0] & !a[1] & a[2] & !a[3] & a[4];
        d[22] = !a[0] & a[1] & a[2] & !a[3] & a[4];
        d[23] = a[0] & a[1] & a[2] & !a[3] & a[4];
        d[24] = !a[0] & !a[1] & !a[2] & a[3] & a[4];
        d[25] = a[0] & !a[1] & !a[2] & a[3] & a[4];
        d[26] = !a[0] & a[1] & !a[2] & a[3] & a[4];
        d[27] = a[0] & a[1] & !a[2] & a[3] & a[4]; 
        d[28] = !a[0] & !a[1] & a[2] & a[3] & a[4];
        d[29] = a[0] & !a[1] & a[2] & a[3] & a[4];
        d[30] = !a[0] & a[1] & a[2] & a[3] & a[4];
        d[31] = a[0] & a[1] & a[2] & a[3] & a[4];
      end
    else d = 32'b00000000000000000000000000000000;
  end
endmodule


* /home/inderjitsingh/eSim-2.3/library/SubcircuitLibrary/8_bit_SRAM_sym/8_bit_SRAM_sym.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 12:41:17 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad10_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad11_ 1_bit_SRAM_isd		
X2  Net-_U1-Pad3_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad12_ 1_bit_SRAM_isd		
X3  Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad13_ 1_bit_SRAM_isd		
X4  Net-_U1-Pad5_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad14_ 1_bit_SRAM_isd		
X5  Net-_U1-Pad6_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad15_ 1_bit_SRAM_isd		
X6  Net-_U1-Pad7_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad16_ 1_bit_SRAM_isd		
X7  Net-_U1-Pad8_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad17_ 1_bit_SRAM_isd		
X8  Net-_U1-Pad9_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad18_ 1_bit_SRAM_isd		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad18_ PORT		

.end

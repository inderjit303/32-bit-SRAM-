* /home/inderjitsingh/eSim-2.3/library/SubcircuitLibrary/1bit_sram_sym/1bit_sram_sym.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 02:00:37 AM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ idata_writer_cktsd		
U4  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U4-Pad3_ Net-_U4-Pad4_ dac_bridge_2		
X1  Net-_U4-Pad3_ Net-_U2-Pad1_ Net-_SC1-Pad2_ Net-_U4-Pad4_ 6t_isramsd		
SC2  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__nfet_01v8		
SC3  Net-_SC2-Pad3_ Net-_SC3-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC4  Net-_SC1-Pad1_ Net-_SC3-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
v1  Net-_SC1-Pad3_ GND DC		
SC6  Net-_SC5-Pad1_ Net-_SC1-Pad1_ GND GND sky130_fd_pr__nfet_01v8		
SC5  Net-_SC5-Pad1_ Net-_SC1-Pad1_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_SC3-Pad2_ Net-_SC5-Pad1_ PORT		

.end
